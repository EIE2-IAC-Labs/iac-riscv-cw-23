module 2flipflop (
    input logic         RegWriteD
    input logic         ResultSrcD
    input logic         MemWriteD
    input logic         JumpD
    input logic         BranchD
    input logic         ALUContrlD
    input logic         ALUSrcD
    input logic         ImmSrcD
    input logic         RD1
    input logic         RD2
    input logic         PCD
    input logic         RdD
    input logic         ImmExtD
    input logic         PCPlus4D
    output logic         RegWriteE
    output logic         ResultSrcE
    output logic         MemWriteE
    output logic         JumpE
    output logic         BranchE
    output logic         ALUContrlE
    output logic         ALUSrcE
    output logic         ImmSrcE
    output logic         RD1E
    output logic         RD2E
    output logic         PCE
    output logic         RdE
    output logic         ImmExtE
    output logic         PCPlus4E
)

