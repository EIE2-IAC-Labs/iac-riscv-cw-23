module DataMemory #(
    parameter ADDRESS_WIDTH = 32,
              DATA_WIDTH = 32
)(
    input logic             clk,
    input logic             WE,
    input logic 

)

endmodule