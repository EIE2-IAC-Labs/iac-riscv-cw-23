module 4flipflop (
    input logic         
);

endmodule