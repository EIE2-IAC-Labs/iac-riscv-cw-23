module 3flipflop(
    input logic         clk;
    input logic         ALUOut;
    input logic         
);

endmodule